module
add()

assign add(wire1, wire2, adder);

endmodule
